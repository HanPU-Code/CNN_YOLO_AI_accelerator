module conv_layer 
(
    input   wire                         clk_i,
    input   wire                         rst_n,
    input   wire  [27 * 8 - 1:0]         in_data,
    output  reg   [64 * 16 - 1:0]        out_data   // 원래 64bit
);

    wire [64:0]  c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15;

    sys_array #(       
        .K0       (72'h01_01_01_01_01_01_01_01_01),
        .K1       (72'h01_01_01_01_01_01_01_01_01),
        .K2       (72'h01_01_01_01_01_01_01_01_01),
        .K3       (72'h01_01_01_01_01_01_01_01_01),
        .K4       (72'h01_01_01_01_01_01_01_01_01),
        .K5       (72'h01_01_01_01_01_01_01_01_01),
        .K6       (72'h01_01_01_01_01_01_01_01_01),
        .K7       (72'h01_01_01_01_01_01_01_01_01),
        .K8       (72'h01_01_01_01_01_01_01_01_01),
        .K9       (72'h01_01_01_01_01_01_01_01_01),
        .K10      (72'h01_01_01_01_01_01_01_01_01),
        .K11      (72'h01_01_01_01_01_01_01_01_01),
        .K12      (72'h01_01_01_01_01_01_01_01_01),
        .K13      (72'h01_01_01_01_01_01_01_01_01),
        .K14      (72'h01_01_01_01_01_01_01_01_01),
        .K15      (72'h01_01_01_01_01_01_01_01_01)
    )
    sys_array_0 (
            .clk_i          (clk_i),
            .rst_n          (rst_n),

            .a0             (in_data),

            .c0             (c0 ),
            .c1             (c1 ),
            .c2             (c2 ),
            .c3             (c3 ),
            .c4             (c4 ),
            .c5             (c5 ),
            .c6             (c6 ),
            .c7             (c7 ),
            .c8             (c8 ),
            .c9             (c9 ),
            .c10            (c10),
            .c11            (c11),
            .c12            (c12),
            .c13            (c13),
            .c14            (c14),
            .c15            (c15)
    );

    always @(posedge clk_i) begin
        if (!rst_n) begin
            out_data <= 0;
        end
        else begin
            out_data <= {c0, c1, c2, c3,
                         c4, c5, c6, c7,
                         c8, c9, c10, c11,
                         c12, c13, c14, c15};
        end
    end

endmodule