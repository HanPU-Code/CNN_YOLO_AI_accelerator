`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/08/14 10:20:21
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
input   wire        clk_i,
input   wire        rst_n,
output  wire        done_o
);

conv_layer conv_layer_0 
(
    .clk_i       (clk_i),
    .rst_n       (rst_n),
    .in_data     (),
    .c           ()
);
endmodule
